module alu_tb();  
  reg zx, zy, nx, ny, f, no;
  reg[7:0] X;
  reg[7:0] Y;
  wire[7:0] O;
  alu alu1 (zx, nx, zy, ny, f, no, X, Y, O);

  initial begin
  $display("zx nx zy ny f no X Y O");
  zx=0; nx=0; zy=1; ny=0; f=1; no=0; X=20; Y=15; #20;
  $display("X:%d Y:%d -> X -> output -> %d", X, Y, O);
  #10;
  zx=1; nx=0; zy=0; ny=0; f=1; no=0; X=20; Y=15; #20;
  $display("X:%d Y:%d -> Y -> output -> %d", X, Y, O);
  #10;
  zx=0; nx=0; zy=0; ny=0; f=0; no=0; X=16; Y=17; #20;
  $display("X:%d Y:%d -> X & Y -> output -> %d", X, Y, O);
  #10;
  zx=0; nx=1; zy=0; ny=1; f=0; no=1; X=16; Y=8; #20;
  $display("X:%d Y:%d -> X | Y -> output -> %d", X, Y, O);
  #10;
  zx=0; nx=1; zy=1; ny=0; f=1; no=0; X=1; Y=15; #20;
  $display("X:%d Y:%d -> ~X -> output -> %d", X, Y, O);
  #10;
  zx=0; nx=1; zy=1; ny=0; f=1; no=0; X=13; Y=255; #20;
  $display("X:%d Y:%d -> ~Y -> output -> %d", X, Y, O);
  #10;
  zx=0; nx=0; zy=0; ny=0; f=1; no=0; X=20; Y=15; #20;
  $display("X:%d Y:%d -> X + Y -> output -> %d", X, Y, O);
  #10;
  zx=0; nx=1; zy=0; ny=0; f=1; no=1; X=20; Y=15; #20;
  $display("X:%d Y:%d -> X - Y -> output -> %d", X, Y, O);
  #10;
  zx=0; nx=0; zy=0; ny=1; f=1; no=1; X=20; Y=15; #20;
  $display("X:%d Y:%d -> Y - X -> output -> %d", X, Y, O);
  #10;
  zx=1; nx=0; zy=1; ny=0; f=1; no=0; X=20; Y=15; #20;
  $display("X:%d Y:%d -> 0 -> output -> %d", X, Y, O);
  #10;
  zx=1; nx=1; zy=1; ny=0; f=1; no=0; X=20; Y=15; #20;
  $display("X:%d Y:%d -> -1 -> output -> %d", X, Y, O);
  #10;
  zx=1; nx=1; zy=1; ny=1; f=1; no=1; X=20; Y=15; #20;
  $display("X:%d Y:%d -> 1 -> output -> %d", X, Y, O);
  #10;
  zx=0; nx=0; zy=1; ny=1; f=1; no=1; X=20; Y=15; #20;
  $display("X:%d Y:%d -> -X -> output -> %d", X, Y, O);
  #10;
  zx=1; nx=1; zy=0; ny=0; f=1; no=1; X=20; Y=15; #20;
  $display("X:%d Y:%d -> -Y -> output -> %d", X, Y, O);
  #10;
  zx=0; nx=1; zy=1; ny=1; f=1; no=1; X=20; Y=15; #20;
  $display("X:%d Y:%d -> X + 1 -> output -> %d", X, Y, O);
  #10;
  zx=1; nx=1; zy=0; ny=1; f=1; no=1; X=20; Y=15; #20;
  $display("X:%d Y:%d -> Y + 1 -> output -> %d", X, Y, O);
  #10;
  zx=0; nx=0; zy=1; ny=1; f=1; no=0; X=20; Y=15; #20;
  $display("X:%d Y:%d -> X - 1 -> output -> %d", X, Y, O);
  #10;
  zx=1; nx=1; zy=0; ny=0; f=1; no=0; X=20; Y=15; #20;
  $display("X:%d Y:%d -> Y - 1 -> output -> %d", X, Y, O);
  #10;
  end
endmodule // test
